magic
tech sky130A
timestamp 1726400396
<< nwell >>
rect -880 3240 -794 3253
rect -880 3079 -538 3240
rect -470 2773 -385 2776
rect -470 2772 -376 2773
rect -470 2690 -181 2772
rect -469 2588 -181 2690
rect -467 2526 -181 2588
rect 49 2284 510 2522
rect 49 2276 338 2284
rect 244 2275 338 2276
rect 253 2272 338 2275
rect -973 2048 -631 2209
rect -717 2035 -631 2048
rect -173 245 7 246
rect -173 183 2 245
rect 240 217 288 246
rect -173 9 0 183
rect -173 8 -1 9
<< nmos >>
rect -714 2979 -699 3021
rect 170 2583 209 2633
rect -341 2415 -302 2465
rect -812 2267 -797 2309
<< pmos >>
rect -714 3099 -699 3178
rect -340 2606 -301 2675
rect 169 2373 208 2442
rect -812 2110 -797 2189
<< ndiff >>
rect -774 3006 -714 3021
rect -774 2986 -754 3006
rect -734 2986 -714 3006
rect -774 2979 -714 2986
rect -699 3011 -644 3021
rect -699 2991 -671 3011
rect -651 2991 -644 3011
rect -699 2986 -644 2991
rect -699 2979 -674 2986
rect 80 2633 125 2636
rect 80 2626 170 2633
rect 80 2598 90 2626
rect 119 2598 170 2626
rect 80 2583 170 2598
rect 209 2624 308 2633
rect 209 2596 266 2624
rect 295 2596 308 2624
rect 209 2583 308 2596
rect -440 2452 -341 2465
rect -440 2424 -427 2452
rect -398 2424 -341 2452
rect -440 2415 -341 2424
rect -302 2450 -212 2465
rect -302 2422 -251 2450
rect -222 2422 -212 2450
rect -302 2415 -212 2422
rect -257 2412 -212 2415
rect -837 2302 -812 2309
rect -867 2297 -812 2302
rect -867 2277 -860 2297
rect -840 2277 -812 2297
rect -867 2267 -812 2277
rect -797 2302 -737 2309
rect -797 2282 -777 2302
rect -757 2282 -737 2302
rect -797 2267 -737 2282
<< pdiff >>
rect -775 3205 -598 3222
rect -688 3178 -644 3205
rect -774 3167 -714 3178
rect -774 3147 -754 3167
rect -734 3147 -714 3167
rect -774 3129 -714 3147
rect -774 3109 -754 3129
rect -734 3109 -714 3129
rect -774 3099 -714 3109
rect -699 3167 -644 3178
rect -699 3147 -679 3167
rect -659 3147 -644 3167
rect -699 3129 -644 3147
rect -699 3109 -679 3129
rect -659 3109 -644 3129
rect -699 3099 -644 3109
rect -451 2644 -340 2675
rect -451 2616 -427 2644
rect -398 2616 -340 2644
rect -451 2606 -340 2616
rect -301 2640 -204 2675
rect -301 2612 -248 2640
rect -219 2612 -204 2640
rect -301 2606 -204 2612
rect 72 2436 169 2442
rect 72 2408 87 2436
rect 116 2408 169 2436
rect 72 2373 169 2408
rect 208 2432 446 2442
rect 208 2404 266 2432
rect 295 2404 446 2432
rect 208 2375 446 2404
rect 208 2373 319 2375
rect -867 2179 -812 2189
rect -867 2159 -852 2179
rect -832 2159 -812 2179
rect -867 2141 -812 2159
rect -867 2121 -852 2141
rect -832 2121 -812 2141
rect -867 2110 -812 2121
rect -797 2179 -737 2189
rect -797 2159 -777 2179
rect -757 2159 -737 2179
rect -797 2141 -737 2159
rect -797 2121 -777 2141
rect -757 2121 -737 2141
rect -797 2110 -737 2121
rect -867 2083 -823 2110
rect -913 2066 -736 2083
rect -109 99 18 166
<< ndiffc >>
rect -754 2986 -734 3006
rect -671 2991 -651 3011
rect 90 2598 119 2626
rect 266 2596 295 2624
rect -427 2424 -398 2452
rect -251 2422 -222 2450
rect -860 2277 -840 2297
rect -777 2282 -757 2302
<< pdiffc >>
rect -754 3147 -734 3167
rect -754 3109 -734 3129
rect -679 3147 -659 3167
rect -679 3109 -659 3129
rect -427 2616 -398 2644
rect -248 2612 -219 2640
rect 87 2408 116 2436
rect 266 2404 295 2432
rect -852 2159 -832 2179
rect -852 2121 -832 2141
rect -777 2159 -757 2179
rect -777 2121 -757 2141
<< psubdiff >>
rect -613 3006 -558 3023
rect -613 2986 -595 3006
rect -575 2986 -558 3006
rect -613 2979 -558 2986
rect -953 2302 -898 2309
rect -953 2282 -936 2302
rect -916 2282 -898 2302
rect -953 2265 -898 2282
<< nsubdiff >>
rect -852 3202 -824 3230
rect -612 3166 -557 3177
rect -612 3108 -591 3166
rect -571 3108 -557 3166
rect -612 3098 -557 3108
rect -954 2180 -899 2190
rect -954 2122 -940 2180
rect -920 2122 -899 2180
rect -954 2111 -899 2122
rect -687 2058 -659 2086
<< psubdiffcont >>
rect -595 2986 -575 3006
rect -936 2282 -916 2302
<< nsubdiffcont >>
rect -591 3108 -571 3166
rect -940 2122 -920 2180
<< poly >>
rect -714 3178 -699 3191
rect -714 3071 -699 3099
rect -714 3062 -673 3071
rect -714 3045 -699 3062
rect -682 3045 -673 3062
rect -714 3032 -673 3045
rect -714 3021 -699 3032
rect -714 2966 -699 2979
rect -350 2741 -333 2746
rect 170 2743 209 2751
rect -350 2733 -291 2741
rect -350 2705 -333 2733
rect -304 2705 -291 2733
rect -349 2696 -291 2705
rect 170 2715 175 2743
rect 204 2715 209 2743
rect -340 2675 -301 2696
rect 170 2633 209 2715
rect -340 2559 -301 2606
rect 170 2563 209 2583
rect -341 2465 -302 2485
rect 169 2442 208 2489
rect -341 2333 -302 2415
rect 169 2352 208 2373
rect -812 2309 -797 2322
rect -341 2305 -336 2333
rect -307 2305 -302 2333
rect 159 2343 217 2352
rect 159 2315 172 2343
rect 201 2315 218 2343
rect 159 2307 218 2315
rect -341 2297 -302 2305
rect 201 2302 218 2307
rect -812 2256 -797 2267
rect -838 2243 -797 2256
rect -838 2226 -829 2243
rect -812 2226 -797 2243
rect -838 2217 -797 2226
rect -812 2189 -797 2217
rect -812 2097 -797 2110
rect 145 451 149 458
<< polycont >>
rect -699 3045 -682 3062
rect -333 2705 -304 2733
rect 175 2715 204 2743
rect -336 2305 -307 2333
rect 172 2315 201 2343
rect -829 2226 -812 2243
<< locali >>
rect -775 3205 -679 3222
rect -688 3201 -679 3205
rect -658 3205 -598 3222
rect -658 3201 -644 3205
rect -688 3177 -644 3201
rect -688 3174 -562 3177
rect -764 3167 -724 3174
rect -764 3147 -754 3167
rect -734 3147 -724 3167
rect -764 3129 -724 3147
rect -764 3109 -754 3129
rect -734 3109 -724 3129
rect -764 3104 -724 3109
rect -689 3167 -562 3174
rect -689 3147 -679 3167
rect -659 3166 -562 3167
rect -659 3147 -591 3166
rect -689 3129 -591 3147
rect -689 3109 -679 3129
rect -659 3109 -591 3129
rect -689 3108 -591 3109
rect -571 3108 -562 3166
rect -689 3104 -562 3108
rect -764 3068 -744 3104
rect -1008 3060 -744 3068
rect -1008 3040 -998 3060
rect -978 3040 -744 3060
rect -1008 3039 -744 3040
rect -707 3064 -543 3067
rect -707 3062 -565 3064
rect -707 3045 -699 3062
rect -682 3047 -565 3062
rect -548 3047 -543 3064
rect -682 3045 -543 3047
rect -707 3039 -543 3045
rect -1008 3038 -972 3039
rect -764 3016 -744 3039
rect -764 3006 -724 3016
rect -764 2986 -754 3006
rect -734 2986 -724 3006
rect -764 2979 -724 2986
rect -689 3011 -564 3016
rect -689 2991 -671 3011
rect -651 3006 -564 3011
rect -651 2991 -595 3006
rect -689 2986 -595 2991
rect -575 2986 -564 3006
rect -689 2979 -564 2986
rect -689 2953 -644 2979
rect -785 2931 -783 2952
rect -689 2932 -676 2953
rect -655 2932 -644 2953
rect -689 2931 -644 2932
rect -785 2897 -762 2931
rect -847 2896 -762 2897
rect -847 2875 -827 2896
rect -806 2875 -762 2896
rect -847 2872 -762 2875
rect 154 2848 215 2849
rect -292 2847 -114 2848
rect -42 2847 215 2848
rect -343 2820 215 2847
rect 1417 2822 1438 2826
rect 318 2820 1438 2822
rect -343 2815 1438 2820
rect -343 2807 240 2815
rect -343 2806 -114 2807
rect -91 2806 240 2807
rect -343 2756 -292 2806
rect -91 2805 -44 2806
rect 154 2794 240 2806
rect 261 2814 1438 2815
rect 261 2794 1445 2814
rect 154 2783 1445 2794
rect -350 2733 -291 2756
rect 154 2751 215 2783
rect 318 2774 1445 2783
rect 154 2749 228 2751
rect -350 2705 -333 2733
rect -304 2705 -291 2733
rect -349 2696 -291 2705
rect 159 2743 228 2749
rect 159 2715 175 2743
rect 204 2715 228 2743
rect 159 2702 228 2715
rect -435 2656 -391 2690
rect -435 2644 -390 2656
rect -435 2616 -427 2644
rect -398 2616 -390 2644
rect -1283 2580 -821 2593
rect -1283 2559 -852 2580
rect -831 2559 -821 2580
rect -435 2560 -390 2616
rect -1283 2545 -821 2559
rect -558 2552 -390 2560
rect -1283 493 -1221 2545
rect -558 2532 -517 2552
rect -497 2532 -390 2552
rect -558 2527 -390 2532
rect -558 2521 -461 2527
rect -435 2452 -390 2527
rect -257 2645 -213 2649
rect -257 2640 -212 2645
rect -257 2612 -248 2640
rect -219 2612 -212 2640
rect -257 2559 -212 2612
rect 80 2626 125 2636
rect 261 2631 303 2657
rect 80 2598 90 2626
rect 119 2598 125 2626
rect -257 2526 -186 2559
rect -260 2524 -184 2526
rect -260 2496 -225 2524
rect -196 2522 -184 2524
rect 80 2522 125 2598
rect -196 2496 -114 2522
rect -260 2494 -114 2496
rect 49 2521 125 2522
rect -260 2493 -121 2494
rect 49 2493 62 2521
rect 91 2493 125 2521
rect -435 2424 -427 2452
rect -398 2424 -390 2452
rect -435 2417 -390 2424
rect -257 2450 -212 2493
rect 54 2489 125 2493
rect -257 2422 -251 2450
rect -222 2422 -212 2450
rect -435 2391 -393 2417
rect -257 2412 -212 2422
rect 80 2436 125 2489
rect 80 2408 87 2436
rect 116 2408 125 2436
rect 80 2403 125 2408
rect 81 2399 125 2403
rect 258 2624 303 2631
rect 258 2596 266 2624
rect 295 2596 303 2624
rect 258 2566 303 2596
rect 258 2538 272 2566
rect 301 2538 303 2566
rect 258 2521 303 2538
rect 258 2488 330 2521
rect 258 2432 303 2488
rect 258 2404 266 2432
rect 295 2404 303 2432
rect 258 2392 303 2404
rect 259 2358 303 2392
rect -867 2356 -847 2357
rect -867 2335 -856 2356
rect -835 2335 -822 2356
rect -867 2309 -822 2335
rect -360 2333 -291 2346
rect -947 2302 -822 2309
rect -947 2282 -936 2302
rect -916 2297 -822 2302
rect -916 2282 -860 2297
rect -947 2277 -860 2282
rect -840 2277 -822 2297
rect -947 2272 -822 2277
rect -787 2302 -747 2309
rect -787 2282 -777 2302
rect -757 2282 -747 2302
rect -360 2305 -336 2333
rect -307 2305 -291 2333
rect -360 2297 -291 2305
rect 159 2343 217 2352
rect 159 2315 172 2343
rect 201 2315 218 2343
rect 159 2302 218 2315
rect -787 2272 -747 2282
rect -767 2256 -747 2272
rect -345 2256 -313 2297
rect 157 2276 217 2302
rect -767 2250 -563 2256
rect -838 2247 -804 2249
rect -1009 2245 -804 2247
rect -1009 2225 -1003 2245
rect -983 2243 -804 2245
rect -983 2226 -829 2243
rect -812 2226 -804 2243
rect -983 2225 -804 2226
rect -1009 2221 -804 2225
rect -767 2230 -589 2250
rect -569 2230 -563 2250
rect -767 2225 -563 2230
rect -344 2235 -313 2256
rect 156 2250 206 2276
rect 156 2248 268 2250
rect 156 2235 224 2248
rect -344 2233 -82 2235
rect -43 2233 224 2235
rect -344 2227 224 2233
rect 245 2227 268 2248
rect -344 2225 268 2227
rect -1009 2220 -837 2221
rect -767 2184 -747 2225
rect -344 2213 206 2225
rect -949 2180 -822 2184
rect -949 2122 -940 2180
rect -920 2179 -822 2180
rect -920 2159 -852 2179
rect -832 2159 -822 2179
rect -920 2141 -822 2159
rect -920 2122 -852 2141
rect -949 2121 -852 2122
rect -832 2121 -822 2141
rect -949 2114 -822 2121
rect -787 2179 -747 2184
rect -787 2159 -777 2179
rect -757 2159 -747 2179
rect -787 2141 -747 2159
rect -787 2121 -777 2141
rect -757 2121 -747 2141
rect -122 2171 -94 2213
rect -122 2150 -119 2171
rect -98 2150 -94 2171
rect -122 2134 -94 2150
rect -787 2114 -747 2121
rect -949 2111 -823 2114
rect -867 2087 -823 2111
rect -867 2083 -853 2087
rect -913 2066 -853 2083
rect -832 2083 -823 2087
rect -832 2066 -736 2083
rect 1299 1005 1344 1014
rect 1299 985 1309 1005
rect 1329 985 1344 1005
rect -566 960 935 967
rect -644 952 935 960
rect -644 931 899 952
rect 920 938 935 952
rect 920 935 937 938
rect 920 931 995 935
rect -644 925 995 931
rect -644 904 -622 925
rect -601 921 995 925
rect -601 904 -567 921
rect -644 894 -567 904
rect 1299 792 1344 985
rect 880 788 1010 791
rect 880 771 885 788
rect 902 771 1010 788
rect 880 763 1010 771
rect 1085 784 1345 792
rect 1085 764 1315 784
rect 1335 764 1345 784
rect 1085 763 1345 764
rect 1309 762 1345 763
rect 67 671 178 680
rect 832 672 917 673
rect 67 664 798 671
rect 67 643 84 664
rect 105 651 798 664
rect 819 655 917 672
rect 1120 655 1122 676
rect 819 651 849 655
rect 105 649 849 651
rect 105 643 178 649
rect 67 632 178 643
rect 773 622 802 649
rect 773 621 819 622
rect 1099 621 1122 655
rect 773 620 1184 621
rect 773 605 1143 620
rect 774 599 1143 605
rect 1164 599 1184 620
rect 774 597 1184 599
rect 1099 596 1184 597
rect 122 572 183 573
rect 122 571 379 572
rect 451 571 629 572
rect 122 565 680 571
rect 122 544 297 565
rect 318 558 680 565
rect 318 544 640 558
rect 11 539 640 544
rect 11 518 76 539
rect 97 537 640 539
rect 661 537 680 558
rect 97 531 680 537
rect 97 530 428 531
rect 451 530 680 531
rect 97 518 183 530
rect 381 529 428 530
rect 11 507 183 518
rect -1276 82 -1221 493
rect 105 488 183 507
rect 107 473 183 488
rect 629 480 680 530
rect 107 469 122 473
rect 149 468 160 473
rect 628 469 687 480
rect 145 451 149 458
rect 1417 441 1445 2774
rect 1424 440 1445 441
rect -431 394 -377 402
rect -431 373 -408 394
rect -387 373 -377 394
rect -730 183 -662 186
rect -730 162 -704 183
rect -683 162 -662 183
rect -730 159 -662 162
rect -572 182 -542 191
rect -572 161 -570 182
rect -549 161 -542 182
rect -572 149 -542 161
rect -431 111 -377 373
rect 1142 304 1184 316
rect 798 276 895 284
rect 798 256 834 276
rect 854 256 895 276
rect 521 248 597 250
rect 521 246 533 248
rect 240 245 288 246
rect 240 217 246 245
rect 275 217 288 245
rect 451 220 533 246
rect 562 220 597 248
rect 798 245 895 256
rect 1142 283 1151 304
rect 1172 283 1184 304
rect 451 218 597 220
rect 458 217 597 218
rect -431 95 -388 111
rect -1278 81 -691 82
rect -1278 47 -686 81
rect -431 74 -417 95
rect -396 74 -388 95
rect 1142 80 1184 283
rect -431 69 -388 74
rect -1269 43 -686 47
rect -1269 42 -705 43
rect -809 31 -778 42
rect -809 15 -804 31
rect -783 15 -778 31
rect -432 8 -388 69
rect 120 0 180 26
rect 131 -26 181 0
rect 69 -28 181 -26
rect 69 -49 92 -28
rect 113 -41 181 -28
rect 650 -20 682 31
rect 421 -38 459 -29
rect 421 -41 430 -38
rect 113 -43 380 -41
rect 419 -43 430 -41
rect 113 -49 430 -43
rect 69 -51 430 -49
rect 131 -59 430 -51
rect 451 -41 459 -38
rect 650 -41 681 -20
rect 451 -59 681 -41
rect 900 -26 1104 -20
rect 900 -46 906 -26
rect 926 -46 1104 -26
rect 900 -51 1104 -46
rect 1174 -31 1346 -29
rect 1174 -51 1320 -31
rect 1340 -51 1346 -31
rect 1174 -56 1346 -51
rect 131 -63 681 -59
rect 1424 -313 1448 440
rect 431 -323 1448 -313
rect 431 -344 435 -323
rect 456 -344 1448 -323
rect 431 -360 1448 -344
rect 1424 -362 1448 -360
<< viali >>
rect -679 3201 -658 3222
rect -998 3040 -978 3060
rect -565 3047 -548 3064
rect -783 2931 -762 2952
rect -676 2932 -655 2953
rect -827 2875 -806 2896
rect 240 2794 261 2815
rect -852 2559 -831 2580
rect -517 2532 -497 2552
rect -225 2496 -196 2524
rect 62 2493 91 2521
rect 272 2538 301 2566
rect -856 2335 -835 2356
rect -1003 2225 -983 2245
rect -589 2230 -569 2250
rect 224 2227 245 2248
rect -119 2150 -98 2171
rect -853 2066 -832 2087
rect 1309 985 1329 1005
rect 899 931 920 952
rect -622 904 -601 925
rect 885 771 902 788
rect 1315 764 1335 784
rect 84 643 105 664
rect 798 651 819 672
rect 1099 655 1120 676
rect 1143 599 1164 620
rect 297 544 318 565
rect 76 518 97 539
rect 640 537 661 558
rect -408 373 -387 394
rect -704 162 -683 183
rect -570 161 -549 182
rect 36 262 65 290
rect 834 256 854 276
rect 246 217 275 245
rect 533 220 562 248
rect 1151 283 1172 304
rect -417 74 -396 95
rect -804 10 -783 31
rect 92 -49 113 -28
rect 430 -59 451 -38
rect 906 -46 926 -26
rect 1320 -51 1340 -31
rect 435 -344 456 -323
<< metal1 >>
rect -1045 3242 -582 3243
rect -1045 3222 -579 3242
rect -1045 3201 -679 3222
rect -658 3201 -579 3222
rect -1045 3193 -579 3201
rect -1045 3191 -582 3193
rect -1045 3190 -1024 3191
rect -1045 2106 -1026 3190
rect -849 3179 -582 3191
rect -849 3178 -644 3179
rect -599 3178 -582 3179
rect -1007 3060 -973 3066
rect -1007 3040 -998 3060
rect -978 3040 -973 3060
rect -573 3064 -524 3067
rect -573 3047 -565 3064
rect -548 3056 -524 3064
rect -548 3047 -83 3056
rect -573 3043 -83 3047
rect -542 3040 -83 3043
rect -1007 3038 -973 3040
rect -1011 2245 -972 3038
rect -689 2979 -674 2986
rect -776 2974 -574 2979
rect -792 2961 -574 2974
rect -113 2971 -83 3040
rect -792 2960 -598 2961
rect -790 2953 -598 2960
rect -790 2952 -676 2953
rect -790 2931 -783 2952
rect -762 2932 -676 2952
rect -655 2932 -598 2953
rect -762 2931 -598 2932
rect -790 2919 -598 2931
rect -112 2913 -85 2971
rect -849 2896 -797 2902
rect -849 2885 -827 2896
rect -865 2875 -827 2885
rect -806 2875 -797 2896
rect -865 2872 -797 2875
rect -865 2850 -821 2872
rect -860 2580 -821 2850
rect -113 2847 -83 2913
rect -860 2559 -852 2580
rect -831 2559 -821 2580
rect -860 2372 -821 2559
rect -558 2552 -449 2560
rect -558 2532 -517 2552
rect -497 2532 -449 2552
rect -865 2356 -823 2372
rect -865 2335 -856 2356
rect -835 2353 -823 2356
rect -835 2335 -824 2353
rect -865 2323 -824 2335
rect -865 2310 -822 2323
rect -856 2309 -822 2310
rect -837 2302 -822 2309
rect -558 2258 -449 2532
rect -258 2526 -185 2527
rect -259 2524 -184 2526
rect -259 2496 -225 2524
rect -196 2522 -184 2524
rect -114 2522 -91 2847
rect 207 2815 270 2820
rect 207 2794 240 2815
rect 261 2794 270 2815
rect 207 2784 270 2794
rect 207 2774 261 2784
rect 170 2760 261 2774
rect 170 2706 207 2760
rect 260 2568 306 2569
rect 260 2567 324 2568
rect 260 2566 341 2567
rect 260 2538 272 2566
rect 301 2544 1345 2566
rect 301 2538 341 2544
rect 260 2535 341 2538
rect 260 2534 324 2535
rect 49 2522 98 2525
rect 1198 2522 1345 2544
rect -196 2521 98 2522
rect -196 2496 62 2521
rect -259 2494 62 2496
rect -259 2491 -122 2494
rect -91 2493 62 2494
rect 91 2493 98 2521
rect 59 2490 95 2493
rect -1011 2225 -1003 2245
rect -983 2225 -972 2245
rect -1011 2223 -972 2225
rect -1010 2221 -972 2223
rect -593 2250 -449 2258
rect -593 2230 -589 2250
rect -569 2230 -449 2250
rect -593 2213 -449 2230
rect 206 2262 251 2271
rect 206 2248 339 2262
rect 206 2227 224 2248
rect 245 2244 339 2248
rect 245 2227 342 2244
rect 206 2223 342 2227
rect -126 2174 -109 2176
rect 273 2174 342 2223
rect -126 2171 342 2174
rect -126 2150 -119 2171
rect -98 2150 342 2171
rect -126 2147 342 2150
rect -1082 2104 -1026 2106
rect -929 2109 -912 2110
rect -867 2109 -662 2110
rect -929 2106 -662 2109
rect -929 2104 -592 2106
rect -1148 2087 -592 2104
rect -1148 2066 -853 2087
rect -832 2070 -592 2087
rect -832 2066 -579 2070
rect -1148 2052 -579 2066
rect -929 2045 -579 2052
rect -686 2033 -579 2045
rect -647 925 -579 2033
rect -647 904 -622 925
rect -601 921 -579 925
rect -601 904 -569 921
rect -647 902 -569 904
rect -645 610 -569 902
rect -402 687 99 688
rect -402 686 107 687
rect -402 667 110 686
rect -437 664 110 667
rect -437 643 84 664
rect 105 643 110 664
rect -437 625 110 643
rect -437 624 107 625
rect -644 357 -571 610
rect -437 402 -378 624
rect 273 565 342 2147
rect 1308 1345 1341 2522
rect 1315 1258 1341 1345
rect 1315 1227 1350 1258
rect 1315 1164 1345 1227
rect 886 1010 920 1011
rect 886 1007 1250 1010
rect 886 990 1285 1007
rect 886 967 920 990
rect 886 952 922 967
rect 886 931 899 952
rect 920 931 922 952
rect 886 907 922 931
rect 1249 935 1285 990
rect 1300 1005 1345 1164
rect 1300 985 1309 1005
rect 1329 985 1345 1005
rect 1300 981 1345 985
rect 1249 918 1382 935
rect 1282 912 1382 918
rect 861 788 910 791
rect 861 780 885 788
rect 420 771 885 780
rect 902 771 910 788
rect 420 767 910 771
rect 1310 784 1344 790
rect 420 764 879 767
rect 1310 764 1315 784
rect 1335 764 1344 784
rect 420 695 450 764
rect 1310 762 1344 764
rect 422 637 449 695
rect 1072 676 1096 695
rect 1130 685 1135 699
rect 775 675 934 676
rect 775 672 917 675
rect 775 651 798 672
rect 819 655 917 672
rect 819 651 934 655
rect 775 641 934 651
rect 420 571 450 637
rect 1130 629 1186 685
rect 1134 620 1186 629
rect 1134 599 1143 620
rect 1164 599 1186 620
rect -302 544 -253 546
rect 273 544 297 565
rect 318 544 342 565
rect -302 539 130 544
rect -302 518 76 539
rect 97 518 130 539
rect 273 536 342 544
rect -302 506 130 518
rect -302 501 166 506
rect -302 487 167 501
rect -302 484 121 487
rect -437 394 -370 402
rect -437 373 -408 394
rect -387 373 -370 394
rect -437 362 -370 373
rect -644 352 -633 357
rect -628 352 -571 357
rect -644 302 -571 352
rect -302 187 -253 484
rect 106 483 121 484
rect 31 292 77 293
rect 13 290 77 292
rect 13 262 36 290
rect 65 262 77 290
rect 13 258 77 262
rect 239 246 288 249
rect 428 246 451 571
rect 626 558 684 565
rect 626 537 640 558
rect 661 537 684 558
rect 626 419 684 537
rect 1134 304 1186 599
rect 786 276 895 284
rect 786 256 834 276
rect 854 256 895 276
rect 522 250 595 251
rect 521 248 596 250
rect 521 246 533 248
rect 239 245 533 246
rect 239 217 246 245
rect 275 220 533 245
rect 562 220 596 248
rect 275 218 596 220
rect 275 217 428 218
rect 242 214 278 217
rect 459 215 596 218
rect -879 183 -658 187
rect -879 162 -704 183
rect -683 162 -658 183
rect -879 158 -658 162
rect -584 186 -253 187
rect -584 182 -257 186
rect -584 161 -570 182
rect -549 161 -257 182
rect -879 -5 -838 158
rect -584 154 -257 161
rect -542 101 -500 103
rect -542 95 -388 101
rect -542 74 -417 95
rect -396 74 -388 95
rect -754 53 -733 74
rect -506 62 -388 74
rect -811 31 -776 36
rect -811 19 -804 31
rect -810 10 -804 19
rect -783 27 -776 31
rect -432 27 -388 62
rect -783 10 -392 27
rect -810 5 -392 10
rect -879 -13 -837 -5
rect -368 -13 -9 -5
rect -879 -14 -9 -13
rect 86 -14 131 -5
rect -879 -28 131 -14
rect -879 -32 92 -28
rect 55 -49 92 -32
rect 113 -49 131 -28
rect 786 -18 895 256
rect 1134 283 1151 304
rect 1172 283 1186 304
rect 1134 80 1186 283
rect 786 -26 930 -18
rect 55 -53 131 -49
rect 425 -38 457 -32
rect 425 -59 430 -38
rect 451 -59 457 -38
rect 425 -208 457 -59
rect 786 -46 906 -26
rect 926 -46 930 -26
rect 786 -63 930 -46
rect 1309 -31 1348 762
rect 1309 -51 1320 -31
rect 1340 -51 1348 -31
rect 1309 -53 1348 -51
rect 1309 -55 1347 -53
rect 1363 -170 1382 912
rect 425 -323 466 -208
rect 973 -234 999 -170
rect 1363 -172 1419 -170
rect 1266 -224 1485 -172
rect 425 -344 435 -323
rect 456 -344 466 -323
rect 425 -376 466 -344
use assignment2  assignment2_0 ~/Downloads
timestamp 1726379637
transform 1 0 1046 0 1 720
box -171 -77 171 257
use assignment2  assignment2_1
timestamp 1726379637
transform -1 0 1139 0 -1 16
box -171 -77 171 257
use assignment2  assignment2_2
timestamp 1726379637
transform 1 0 -626 0 1 120
box -171 -77 171 257
use tg  tg_0
timestamp 1726386644
transform 0 1 58 -1 0 196
box -279 -59 200 230
use tg  tg_1
timestamp 1726386644
transform 0 -1 748 1 0 300
box -279 -59 200 230
<< labels >>
rlabel viali 44 276 44 276 1 D_in
port 1 n
rlabel viali -559 172 -559 172 1 clk_bar
port 2 n
rlabel viali -696 171 -696 171 1 clock
port 3 n
rlabel viali 1157 292 1157 292 1 GND
port 5 n
rlabel metal1 -633 352 -633 352 1 VDD
port 6 n
rlabel viali 256 236 256 236 1 Q1
port 7 n
rlabel viali 1324 775 1324 775 1 Q1out
port 8 n
rlabel viali 913 -34 913 -34 1 Q1bar_out
port 9 n
rlabel viali 73 2509 73 2509 1 Q1out_bar
port 10 n
rlabel viali -992 3049 -992 3049 1 Q2
port 11 n
<< end >>
