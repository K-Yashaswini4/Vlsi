magic
tech sky130A
timestamp 1726424396
<< nwell >>
rect 1638 1016 1722 1017
rect 1938 1016 2022 1017
rect 1638 858 2282 1016
rect 1638 761 2284 858
rect 1661 760 2284 761
rect 1942 759 2284 760
<< nmos >>
rect 1859 664 1890 706
rect 2020 665 2051 707
<< pmos >>
rect 1859 794 1890 948
rect 2020 793 2051 948
<< ndiff >>
rect 1911 706 2020 707
rect 1781 698 1859 706
rect 1781 678 1787 698
rect 1807 678 1859 698
rect 1781 664 1859 678
rect 1890 703 2020 706
rect 1890 683 1950 703
rect 1970 683 2020 703
rect 1890 665 2020 683
rect 2051 699 2171 707
rect 2051 679 2095 699
rect 2115 679 2171 699
rect 2051 665 2171 679
rect 1890 664 1915 665
rect 1146 342 1198 368
<< pdiff >>
rect 1782 895 1859 948
rect 1782 875 1797 895
rect 1817 875 1859 895
rect 1782 794 1859 875
rect 1890 794 2020 948
rect 1995 793 2020 794
rect 2051 899 2181 948
rect 2051 879 2121 899
rect 2141 879 2181 899
rect 2051 870 2181 879
rect 2051 793 2180 870
<< ndiffc >>
rect 1787 678 1807 698
rect 1950 683 1970 703
rect 2095 679 2115 699
<< pdiffc >>
rect 1797 875 1817 895
rect 2121 879 2141 899
<< psubdiff >>
rect 1681 698 1754 714
rect 1681 678 1708 698
rect 1728 678 1754 698
rect 1681 660 1754 678
<< nsubdiff >>
rect 1669 891 1735 950
rect 1669 871 1690 891
rect 1710 871 1735 891
rect 1669 793 1735 871
<< psubdiffcont >>
rect 1708 678 1728 698
<< nsubdiffcont >>
rect 1690 871 1710 891
<< poly >>
rect 1859 948 1890 970
rect 2020 948 2051 970
rect 1859 748 1890 794
rect 1859 728 1864 748
rect 1884 728 1890 748
rect 1859 706 1890 728
rect 2020 707 2051 793
rect 1859 649 1890 664
rect 2020 649 2051 665
<< polycont >>
rect 1864 728 1884 748
<< locali >>
rect 1780 1054 1830 1062
rect 1780 1034 1794 1054
rect 1814 1034 1830 1054
rect 1780 919 1830 1034
rect 1681 895 1831 919
rect 1681 891 1797 895
rect 1681 871 1690 891
rect 1710 875 1797 891
rect 1817 875 1831 895
rect 1710 871 1831 875
rect 1681 856 1831 871
rect 2106 899 2155 921
rect 2106 879 2121 899
rect 2141 879 2155 899
rect 1841 751 1893 752
rect 2106 751 2155 879
rect 1674 749 1893 751
rect 1674 729 1686 749
rect 1706 748 1893 749
rect 1706 729 1864 748
rect 1674 728 1864 729
rect 1884 728 1893 748
rect 1968 745 2155 751
rect 1674 723 1893 728
rect 1841 722 1893 723
rect 1940 734 2155 745
rect 1699 703 1726 706
rect 1781 703 1812 706
rect 1037 686 1075 699
rect 1037 665 1048 686
rect 1069 665 1075 686
rect 1699 698 1812 703
rect 1940 703 1985 734
rect 1699 678 1708 698
rect 1728 678 1787 698
rect 1807 678 1814 698
rect 1699 673 1814 678
rect 1940 683 1950 703
rect 1970 683 1985 703
rect 1940 677 1985 683
rect 2087 699 2126 707
rect 2087 679 2095 699
rect 2115 679 2126 699
rect 2087 676 2126 679
rect 1699 671 1726 673
rect 1781 670 1814 673
rect 1037 633 1075 665
rect 1786 616 1814 670
rect 2091 662 2124 676
rect 2092 659 2124 662
rect 2092 627 2120 659
rect 1786 596 1790 616
rect 1810 596 1814 616
rect 1786 586 1814 596
rect 2085 620 2121 627
rect 2085 600 2091 620
rect 2111 600 2121 620
rect 2085 589 2121 600
rect 1146 366 1198 368
rect 1146 345 1160 366
rect 1181 345 1198 366
rect 1146 342 1198 345
<< viali >>
rect 1794 1034 1814 1054
rect 1686 729 1706 749
rect 1048 665 1069 686
rect 1790 596 1810 616
rect 2091 600 2111 620
rect 1112 462 1132 482
rect 1160 345 1181 366
<< metal1 >>
rect 1780 1066 1828 1072
rect 1061 1058 1828 1066
rect 1045 1054 1828 1058
rect 1045 1034 1794 1054
rect 1814 1034 1828 1054
rect 1045 879 1072 1034
rect 1780 1031 1828 1034
rect 1040 686 1076 879
rect 1673 749 1715 752
rect 1673 748 1686 749
rect 1348 730 1686 748
rect 1348 723 1398 730
rect 1673 729 1686 730
rect 1706 748 1715 749
rect 1858 748 1891 750
rect 1706 730 1891 748
rect 1706 729 1715 730
rect 1040 665 1048 686
rect 1069 665 1076 686
rect 1040 657 1076 665
rect 1105 482 1139 485
rect 1105 462 1112 482
rect 1132 480 1139 482
rect 1353 480 1383 723
rect 1673 722 1715 729
rect 1858 727 1891 730
rect 1783 617 1827 621
rect 2085 620 2121 627
rect 2085 617 2091 620
rect 1783 616 2091 617
rect 1783 596 1790 616
rect 1810 600 2091 616
rect 2111 600 2121 620
rect 1810 596 2121 600
rect 1783 590 2121 596
rect 1783 589 1827 590
rect 1132 463 1383 480
rect 1132 462 1136 463
rect 1105 457 1136 462
rect 1113 456 1136 457
rect 1891 380 1927 590
rect 2085 589 2121 590
rect 1146 366 1198 368
rect 1146 345 1160 366
rect 1181 345 1198 366
rect 1207 362 1930 380
rect 1146 342 1198 345
use assignment2  assignment2_0
timestamp 1726423755
transform 1 0 1078 0 1 413
box -171 -77 171 257
<< labels >>
rlabel viali 1173 357 1173 357 1 GND
port 1 n
rlabel viali 1059 677 1059 677 1 VDD
port 2 n
rlabel viali 1121 473 1121 473 1 a
port 3 n
rlabel space 1058 468 1058 468 1 abar
port 4 n
rlabel poly 2036 723 2036 723 1 b
port 5 n
<< end >>
