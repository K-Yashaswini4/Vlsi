magic
tech sky130A
timestamp 1726386644
<< nwell >>
rect -50 35 196 230
rect -50 26 197 35
rect -50 -56 200 26
rect 12 -58 200 -56
rect 114 -59 200 -58
<< nmos >>
rect -161 70 -111 109
<< pmos >>
rect 30 71 99 110
<< ndiff >>
rect -164 189 -111 199
rect -164 160 -154 189
rect -126 160 -111 189
rect -164 154 -111 160
rect -161 109 -111 154
rect -161 13 -111 70
rect -161 -16 -152 13
rect -124 -16 -111 13
rect -161 -29 -111 -16
<< pdiff >>
rect 30 192 99 207
rect 30 163 36 192
rect 64 163 99 192
rect 30 110 99 163
rect 30 13 99 71
rect 30 -16 40 13
rect 68 -16 99 13
rect 30 -40 99 -16
<< ndiffc >>
rect -154 160 -126 189
rect -152 -16 -124 13
<< pdiffc >>
rect 36 163 64 192
rect 40 -16 68 13
<< poly >>
rect 120 110 165 120
rect -279 104 -161 109
rect -279 75 -271 104
rect -243 75 -161 104
rect -279 70 -161 75
rect -111 70 -91 109
rect -17 71 30 110
rect 99 107 165 110
rect 99 78 129 107
rect 157 78 165 107
rect 99 71 170 78
rect 120 62 170 71
rect 129 61 170 62
<< polycont >>
rect -271 75 -243 104
rect 129 78 157 107
<< locali >>
rect -50 199 -17 225
rect -164 198 69 199
rect -164 192 73 198
rect -164 189 36 192
rect -164 160 -154 189
rect -126 163 36 189
rect 64 163 73 192
rect -126 160 73 163
rect -164 154 73 160
rect -279 104 -230 120
rect -279 75 -271 104
rect -243 75 -230 104
rect -279 51 -230 75
rect 120 107 170 120
rect 120 78 129 107
rect 157 78 170 107
rect 120 62 170 78
rect 129 61 170 62
rect -159 20 80 21
rect -159 18 114 20
rect -185 13 114 18
rect -185 -16 -152 13
rect -124 -16 40 13
rect 68 -16 114 13
rect -185 -24 114 -16
rect -49 -51 -16 -24
<< end >>
