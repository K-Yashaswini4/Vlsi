* SkyWater PDK
* Simple buffer (inverter-based)

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* Voltage sources:
Vdd vdd gnd DC 1.8
V1 in gnd pulse(0 1.8 0p 200p 100p 1n 2n)

Xnot1 in vdd gnd out1 not1
Xnot2 out1 vdd gnd out not1
.subckt not1 a vdd vss z
xm01	z a	vdd	vdd sky130_fd_pr__pfet_01v8 l=0.15 w=1.1 as=w*l*2 ps=2*(w+2*l) pd=2*(w+2*l)
xm02	z a	vss	vss sky130_fd_pr__nfet_01v8 l=0.15 w=0.4 as=w*l*2 ps=2*(w+2*l) pd=2*(w+2*l)
c3 a vss 0.384f
c2 z vss 0.576f
.ends

* Simulation command:
.tran 1ps 10ns 0 10p
.dc V1 0 1.8 0.01
.control
run
plot in out 
.endc
