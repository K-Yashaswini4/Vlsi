* SkyWater PDK
* Corrected 2-input NOR gate

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* Voltage sources:
Vdd vdd gnd DC 1.8
V1 in1 gnd pulse(0 1.8 0p 200p 100p 1n 2n)
V2 in2 gnd pulse(0 1.8 1n 200p 100p 1n 2n)

Xnor1 in1 in2 vdd gnd out nor

* Corrected NOR gate structure with PMOS in series and NMOS in parallel


.subckt nor a b vdd gnd z
* PMOS transistors in series
xm01	a_bar a	vdd	vdd sky130_fd_pr__pfet_01v8 l=0.15 w=1.1 as=w*l*2 ps=2*(w+2*l) pd=2*(w+2*l)
xm02	a_bar a	gnd	gnd sky130_fd_pr__nfet_01v8 l=0.15 w=0.4 as=w*l*2 ps=2*(w+2*l) pd=2*(w+2*l)
xm03	k a_bar	vdd	vdd sky130_fd_pr__pfet_01v8 l=0.15 w=2.2 as=w*l*2 ps=2*(w+2*l) pd=2*(w+2*l)
xm04	z b	k	k sky130_fd_pr__pfet_01v8 l=0.15 w=2.2 as=w*l*2 ps=2*(w+2*l) pd=2*(w+2*l)
* NMOS transistors in parallel
xm05	z a_bar	gnd	gnd sky130_fd_pr__nfet_01v8 l=0.15 w=0.4 as=w*l*2 ps=2*(w+2*l) pd=2*(w+2*l)
xm06	z b	gnd	gnd sky130_fd_pr__nfet_01v8 l=0.15 w=0.4 as=w*l*2 ps=2*(w+2*l) pd=2*(w+2*l)
* Capacitances for balancing rise/fall times

.ends

* Simulation command:
.tran 1ps 10ns 0 10p
.dc V1 0 1.8 0.01
.dc V2 0 1.8 0.01
.control
run
plot in1 in2 out
.endc
