* SkyWater PDK
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* Voltage sources:
Vdd VDD gnd DC 1.8
V1 in gnd pulse(1.8 1.8 0p 10p 10p 1n 2n)



* Buffer subcircuit
Xnot1 in VDD gnd out not1

* Define subcircuit: Inverter
.subckt not1 A VDD VSS Y2

* Pull-down NMOS transistor
X0 A2 A VSS VSS sky130_fd_pr__nfet_01v8 ad=0.252 pd=2.04 as=0.768847 ps=6.225883 w=0.42 l=0.15
* Pull-up PMOS transistor
X1 A2 A VDD VDD sky130_fd_pr__pfet_01v8 ad=0.474 pd=2.78 as=0.884353 ps=6.260377 w=0.79 l=0.15
* Output stage: Pull-up
X2 Y2 A2 VDD VDD sky130_fd_pr__pfet_01v8 ad=0.432 pd=2.68 as=0.895547 ps=6.339623 w=0.8 l=0.15
* Output stage: Pull-down
X3 Y2 A2 VSS VSS sky130_fd_pr__nfet_01v8 ad=0.2838 pd=2.18 as=0.787153 ps=6.374118 w=0.43 l=0.15

* Parasitic capacitances
C0 Y2 A2 0.040556f
C1 VDD A 0.090563f
C2 A2 A 0.043327f
C3 A2 VDD 0.486332f
C4 Y2 A 2.57e-21
C5 Y2 VDD 0.122326f
C6 Y2 VSS 0.159611f
C7 A2 VSS 0.814371f
C8 A VSS 0.223025f
C9 VDD VSS 2.20592f
.ends

.tran 1ps 100ns 0 10p
*.dc V1 0 1.8 0.01

.control
run
print i(vdd)*1.8
plot i(vdd)*1.8
.endc
