VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO assignment2
  CLASS BLOCK ;
  FOREIGN assignment2 ;
  ORIGIN 1.710 0.800 ;
  SIZE 8.670 BY 3.440 ;
  PIN A
    ANTENNAGATEAREA 0.181500 ;
    PORT
      LAYER li1 ;
        RECT -0.360 0.430 -0.020 0.710 ;
    END
  END A
  PIN Y
    ANTENNAGATEAREA 0.184500 ;
    ANTENNADIFFAREA 0.726000 ;
    PORT
      LAYER li1 ;
        RECT 0.150 1.080 0.550 1.780 ;
        RECT 0.350 0.800 0.550 1.080 ;
        RECT 0.350 0.270 0.800 0.800 ;
        RECT 4.030 0.660 4.520 0.720 ;
        RECT 4.030 0.400 5.100 0.660 ;
        RECT 0.350 0.200 0.550 0.270 ;
        RECT 0.150 -0.170 0.550 0.200 ;
      LAYER met1 ;
        RECT 0.410 0.730 1.200 0.770 ;
        RECT 0.410 0.450 5.100 0.730 ;
        RECT 0.410 0.330 1.200 0.450 ;
        RECT 3.990 0.400 5.100 0.450 ;
    END
  END Y
  PIN VDD
    ANTENNADIFFAREA 2.794700 ;
    PORT
      LAYER nwell ;
        RECT 6.020 2.590 6.960 2.640 ;
        RECT 0.850 2.440 1.710 2.570 ;
        RECT 4.470 2.470 6.960 2.590 ;
        RECT 3.910 2.460 6.960 2.470 ;
        RECT -1.710 0.830 1.710 2.440 ;
        RECT 3.600 2.420 6.960 2.460 ;
        RECT 3.050 1.970 6.960 2.420 ;
        RECT 3.040 1.800 6.960 1.970 ;
        RECT 3.040 0.820 6.860 1.800 ;
        RECT 3.050 0.810 6.860 0.820 ;
      LAYER li1 ;
        RECT -1.110 2.090 0.660 2.260 ;
        RECT 4.110 2.100 5.870 2.270 ;
        RECT -0.650 1.810 -0.210 2.090 ;
        RECT -1.470 1.780 -0.210 1.810 ;
        RECT -1.470 1.080 -0.200 1.780 ;
        RECT 4.470 1.700 4.920 2.100 ;
        RECT 3.390 1.100 4.920 1.700 ;
        RECT 4.470 1.090 4.920 1.100 ;
        RECT 4.470 1.010 4.910 1.090 ;
      LAYER met1 ;
        RECT -1.270 2.460 3.600 2.470 ;
        RECT 3.910 2.460 6.580 2.470 ;
        RECT -1.270 2.210 6.580 2.460 ;
        RECT -1.270 2.020 6.630 2.210 ;
        RECT -1.270 1.830 1.400 2.020 ;
        RECT -1.270 1.820 -1.100 1.830 ;
        RECT -0.650 1.820 1.400 1.830 ;
        RECT 3.600 1.930 6.630 2.020 ;
        RECT 3.600 1.830 6.580 1.930 ;
        RECT 3.600 1.810 4.470 1.830 ;
        RECT 4.920 1.810 6.580 1.830 ;
        RECT 3.600 1.800 3.910 1.810 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 1.021000 ;
    PORT
      LAYER li1 ;
        RECT -1.450 -0.170 -0.200 0.200 ;
        RECT -0.650 -0.450 -0.200 -0.170 ;
        RECT -1.290 -0.650 0.820 -0.450 ;
      LAYER met1 ;
        RECT -1.350 -0.350 1.360 -0.170 ;
        RECT -1.350 -0.630 1.400 -0.350 ;
        RECT -1.350 -0.770 1.360 -0.630 ;
    END
  END VSS
  PIN Y2
    ANTENNADIFFAREA 0.715800 ;
    PORT
      LAYER li1 ;
        RECT 5.240 1.060 5.640 1.760 ;
        RECT 5.390 1.010 5.640 1.060 ;
        RECT 5.440 0.190 5.640 1.010 ;
        RECT 5.240 -0.180 5.640 0.190 ;
    END
  END Y2
  OBS
      LAYER li1 ;
        RECT 4.520 0.170 4.920 0.190 ;
        RECT 3.900 0.150 4.920 0.170 ;
        RECT 3.880 -0.100 4.920 0.150 ;
        RECT 4.520 -0.560 4.920 -0.100 ;
        RECT 4.150 -0.760 6.260 -0.560 ;
      LAYER met1 ;
        RECT 4.520 -0.210 4.920 0.190 ;
        RECT 3.960 -0.800 6.670 -0.210 ;
  END
END assignment2
END LIBRARY

