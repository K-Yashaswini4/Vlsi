magic
tech sky130A
timestamp 1726379637
<< nwell >>
rect 85 244 171 257
rect -171 83 171 244
<< nmos >>
rect -10 -17 5 25
<< pmos >>
rect -10 103 5 182
<< ndiff >>
rect -65 15 -10 25
rect -65 -5 -58 15
rect -38 -5 -10 15
rect -65 -10 -10 -5
rect -35 -17 -10 -10
rect 5 10 65 25
rect 5 -10 25 10
rect 45 -10 65 10
rect 5 -17 65 -10
<< pdiff >>
rect -111 209 66 226
rect -65 182 -21 209
rect -65 171 -10 182
rect -65 151 -50 171
rect -30 151 -10 171
rect -65 133 -10 151
rect -65 113 -50 133
rect -30 113 -10 133
rect -65 103 -10 113
rect 5 171 65 182
rect 5 151 25 171
rect 45 151 65 171
rect 5 133 65 151
rect 5 113 25 133
rect 45 113 65 133
rect 5 103 65 113
<< ndiffc >>
rect -58 -5 -38 15
rect 25 -10 45 10
<< pdiffc >>
rect -50 151 -30 171
rect -50 113 -30 133
rect 25 151 45 171
rect 25 113 45 133
<< psubdiff >>
rect -151 10 -96 27
rect -151 -10 -134 10
rect -114 -10 -96 10
rect -151 -17 -96 -10
<< nsubdiff >>
rect 115 206 143 234
rect -152 170 -97 181
rect -152 112 -138 170
rect -118 112 -97 170
rect -152 102 -97 112
<< psubdiffcont >>
rect -134 -10 -114 10
<< nsubdiffcont >>
rect -138 112 -118 170
<< poly >>
rect -10 182 5 195
rect -10 75 5 103
rect -36 66 5 75
rect -36 49 -27 66
rect -10 49 5 66
rect -36 36 5 49
rect -10 25 5 36
rect -10 -30 5 -17
<< polycont >>
rect -27 49 -10 66
<< locali >>
rect -111 209 -51 226
rect -65 205 -51 209
rect -30 209 66 226
rect -30 205 -21 209
rect -65 181 -21 205
rect -147 178 -21 181
rect -147 171 -20 178
rect -147 170 -50 171
rect -147 112 -138 170
rect -118 151 -50 170
rect -30 151 -20 171
rect -118 133 -20 151
rect -118 113 -50 133
rect -30 113 -20 133
rect -118 112 -20 113
rect -147 108 -20 112
rect 15 171 55 178
rect 15 151 25 171
rect 45 151 55 171
rect 15 133 55 151
rect 15 113 25 133
rect 45 113 55 133
rect 15 108 55 113
rect -36 66 -2 71
rect -36 49 -27 66
rect -10 49 -2 66
rect -36 43 -2 49
rect 35 20 55 108
rect -145 15 -20 20
rect -145 10 -58 15
rect -145 -10 -134 10
rect -114 -5 -58 10
rect -38 -5 -20 15
rect -114 -10 -20 -5
rect -145 -17 -20 -10
rect 15 10 55 20
rect 15 -10 25 10
rect 45 -10 55 10
rect 15 -17 55 -10
rect -65 -43 -20 -17
rect -65 -64 -54 -43
rect -33 -64 -20 -43
rect -65 -65 -20 -64
<< viali >>
rect -51 205 -30 226
rect -54 -64 -33 -43
<< metal1 >>
rect -127 234 140 247
rect -127 226 143 234
rect -127 205 -51 226
rect -30 206 143 226
rect -30 205 140 206
rect -127 183 140 205
rect -127 182 -110 183
rect -65 182 140 183
rect -35 -17 -20 -10
rect -135 -43 84 -17
rect -135 -64 -54 -43
rect -33 -64 84 -43
rect -135 -77 84 -64
<< end >>
