magic
tech sky130A
timestamp 1726080774
<< nwell >>
rect 602 259 696 264
rect 85 244 171 257
rect 447 247 696 259
rect 391 246 696 247
rect -171 83 171 244
rect 360 242 696 246
rect 305 197 696 242
rect 304 180 696 197
rect 304 82 686 180
rect 305 81 686 82
<< nmos >>
rect -10 -17 5 25
rect 502 -21 517 22
<< pmos >>
rect -10 103 5 182
rect 502 101 517 181
<< ndiff >>
rect -65 10 -10 25
rect -65 -10 -50 10
rect -30 -10 -10 10
rect -65 -17 -10 -10
rect 5 10 65 25
rect 5 -10 25 10
rect 45 -10 65 10
rect 5 -17 65 -10
rect 452 4 502 22
rect 452 -16 461 4
rect 481 -16 502 4
rect -65 -45 -20 -17
rect 452 -21 502 -16
rect 517 12 583 22
rect 517 -8 536 12
rect 556 -8 583 12
rect 517 -21 583 -8
rect -129 -65 82 -45
rect 452 -56 492 -21
rect 415 -76 626 -56
<< pdiff >>
rect -111 209 66 226
rect -65 182 -21 209
rect 411 210 587 227
rect -65 171 -10 182
rect -65 151 -50 171
rect -30 151 -10 171
rect -65 133 -10 151
rect -65 113 -50 133
rect -30 113 -10 133
rect -65 103 -10 113
rect 5 171 65 182
rect 447 181 492 210
rect 5 151 25 171
rect 45 151 65 171
rect 5 133 65 151
rect 5 113 25 133
rect 45 113 65 133
rect 5 103 65 113
rect 440 170 502 181
rect 440 150 459 170
rect 479 150 502 170
rect 440 132 502 150
rect 440 112 460 132
rect 480 112 502 132
rect 440 101 502 112
rect 517 169 571 181
rect 517 149 536 169
rect 556 149 571 169
rect 517 131 571 149
rect 517 111 537 131
rect 557 111 571 131
rect 517 101 571 111
<< ndiffc >>
rect -50 -10 -30 10
rect 25 -10 45 10
rect 461 -16 481 4
rect 536 -8 556 12
<< pdiffc >>
rect -50 151 -30 171
rect -50 113 -30 133
rect 25 151 45 171
rect 25 113 45 133
rect 459 150 479 170
rect 460 112 480 132
rect 536 149 556 169
rect 537 111 557 131
<< psubdiff >>
rect -151 10 -96 27
rect -151 -10 -134 10
rect -114 -10 -96 10
rect -151 -17 -96 -10
rect 380 14 424 26
rect 380 -3 397 14
rect 417 -3 424 14
rect 380 -15 424 -3
<< nsubdiff >>
rect 115 206 143 234
rect -152 170 -97 181
rect -152 112 -138 170
rect -118 112 -97 170
rect -152 102 -97 112
rect 635 193 663 221
rect 332 165 387 178
rect 332 117 348 165
rect 384 117 387 165
rect 332 101 387 117
<< psubdiffcont >>
rect -134 -10 -114 10
rect 397 -3 417 14
<< nsubdiffcont >>
rect -138 112 -118 170
rect 348 117 384 165
<< poly >>
rect -10 182 5 195
rect 502 181 517 195
rect -10 75 5 103
rect -36 66 5 75
rect 502 69 517 101
rect -36 49 -27 66
rect -10 49 5 66
rect -36 36 5 49
rect -10 25 5 36
rect 450 61 517 69
rect 450 44 485 61
rect 502 44 517 61
rect 450 30 517 44
rect 502 22 517 30
rect -10 -30 5 -17
rect 502 -34 517 -21
<< polycont >>
rect -27 49 -10 66
rect 485 44 502 61
<< locali >>
rect 411 226 587 227
rect -111 209 -51 226
rect -65 205 -51 209
rect -30 209 66 226
rect 411 210 455 226
rect -30 205 -21 209
rect -65 181 -21 205
rect -147 178 -21 181
rect 447 205 455 210
rect 476 210 587 226
rect 476 205 492 210
rect -147 171 -20 178
rect -147 170 -50 171
rect -147 112 -138 170
rect -118 151 -50 170
rect -30 151 -20 171
rect -118 133 -20 151
rect -118 113 -50 133
rect -30 113 -20 133
rect -118 112 -20 113
rect -147 108 -20 112
rect 15 171 55 178
rect 15 151 25 171
rect 45 151 55 171
rect 447 170 492 205
rect 15 133 55 151
rect 15 113 25 133
rect 45 113 55 133
rect 15 108 55 113
rect 339 165 459 170
rect 339 117 348 165
rect 384 150 459 165
rect 479 150 492 170
rect 384 132 492 150
rect 384 117 460 132
rect 339 112 460 117
rect 480 112 492 132
rect 339 110 492 112
rect 35 80 55 108
rect 447 109 492 110
rect 524 169 564 176
rect 524 149 536 169
rect 556 149 564 169
rect 524 131 564 149
rect 524 111 537 131
rect 557 111 564 131
rect 447 101 491 109
rect 524 106 564 111
rect 539 101 564 106
rect -36 66 -2 71
rect -36 49 -27 66
rect -10 49 -2 66
rect -36 43 -2 49
rect 35 65 80 80
rect 35 44 48 65
rect 69 44 80 65
rect 35 27 80 44
rect 403 69 452 72
rect 403 48 415 69
rect 436 66 452 69
rect 436 61 510 66
rect 436 48 485 61
rect 403 44 485 48
rect 502 44 510 61
rect 403 40 510 44
rect 35 20 55 27
rect -145 10 -20 20
rect -145 -10 -134 10
rect -114 -10 -50 10
rect -30 -10 -20 10
rect -145 -17 -20 -10
rect 15 10 55 20
rect 544 19 564 101
rect 452 17 492 19
rect 390 15 492 17
rect 15 -10 25 10
rect 45 -10 55 10
rect 388 14 492 15
rect 388 -3 397 14
rect 417 4 492 14
rect 417 -3 461 4
rect 388 -10 461 -3
rect 15 -17 55 -10
rect 452 -16 461 -10
rect 481 -16 492 4
rect -65 -43 -20 -17
rect -65 -45 -54 -43
rect -129 -64 -54 -45
rect -33 -45 -20 -43
rect -33 -64 82 -45
rect 452 -54 492 -16
rect 524 12 564 19
rect 524 -8 536 12
rect 556 -8 564 12
rect 524 -18 564 -8
rect 452 -56 462 -54
rect -129 -65 82 -64
rect 415 -75 462 -56
rect 483 -56 492 -54
rect 483 -75 626 -56
rect 415 -76 626 -75
<< viali >>
rect -51 205 -30 226
rect 455 205 476 226
rect 48 44 69 65
rect 415 48 436 69
rect -54 -64 -33 -43
rect 462 -75 483 -54
<< metal1 >>
rect -127 246 360 247
rect 391 246 658 247
rect -127 226 658 246
rect -127 205 -51 226
rect -30 205 455 226
rect 476 221 658 226
rect 476 205 663 221
rect -127 202 663 205
rect -127 183 140 202
rect -127 182 -110 183
rect -65 182 140 183
rect 360 193 663 202
rect 360 183 658 193
rect 360 181 447 183
rect 492 181 658 183
rect 360 180 391 181
rect 41 73 120 77
rect 41 69 510 73
rect 41 65 415 69
rect 41 44 48 65
rect 69 48 415 65
rect 436 48 510 69
rect 69 45 510 48
rect 69 44 120 45
rect 41 33 120 44
rect 399 40 510 45
rect -135 -35 136 -17
rect 452 -21 492 19
rect -135 -43 140 -35
rect -135 -64 -54 -43
rect -33 -63 140 -43
rect 396 -54 667 -21
rect -33 -64 136 -63
rect -135 -77 136 -64
rect 396 -75 462 -54
rect 483 -75 667 -54
rect 396 -80 667 -75
<< labels >>
rlabel locali -36 57 -36 57 7 A
port 1 w
rlabel metal1 -111 217 -111 217 7 VDD
port 3 w
rlabel metal1 -129 -55 -129 -55 7 VSS
port 4 w
rlabel viali 54 56 54 56 3 Y
port 2 e
rlabel locali 478 52 478 52 3 A2
port 6 e
rlabel locali 557 57 557 57 7 Y2
port 7 w
rlabel viali 468 -63 468 -63 1 VSS
<< end >>
