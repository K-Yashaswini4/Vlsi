VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO nor
  CLASS BLOCK ;
  FOREIGN nor ;
  ORIGIN -9.070 -3.360 ;
  SIZE 13.770 BY 7.360 ;
  PIN GND
    ANTENNADIFFAREA 2.358000 ;
    PORT
      LAYER li1 ;
        RECT 16.990 7.030 17.260 7.060 ;
        RECT 17.810 7.030 18.120 7.060 ;
        RECT 16.990 6.980 18.120 7.030 ;
        RECT 16.990 6.730 18.140 6.980 ;
        RECT 20.870 6.760 21.260 7.070 ;
        RECT 16.990 6.710 17.260 6.730 ;
        RECT 17.810 6.700 18.140 6.730 ;
        RECT 17.860 5.860 18.140 6.700 ;
        RECT 20.910 6.620 21.240 6.760 ;
        RECT 20.920 6.590 21.240 6.620 ;
        RECT 20.920 6.270 21.200 6.590 ;
        RECT 20.850 5.890 21.210 6.270 ;
        RECT 9.330 3.960 10.580 4.330 ;
        RECT 10.130 3.680 10.580 3.960 ;
        RECT 9.470 3.480 11.980 3.680 ;
        RECT 11.460 3.420 11.980 3.480 ;
      LAYER met1 ;
        RECT 17.830 6.170 18.270 6.210 ;
        RECT 20.850 6.170 21.210 6.270 ;
        RECT 17.830 5.900 21.210 6.170 ;
        RECT 17.830 5.890 18.270 5.900 ;
        RECT 9.430 3.800 12.140 3.960 ;
        RECT 18.910 3.800 19.270 5.900 ;
        RECT 20.850 5.890 21.210 5.900 ;
        RECT 9.430 3.620 19.300 3.800 ;
        RECT 9.430 3.500 12.180 3.620 ;
        RECT 9.430 3.360 12.140 3.500 ;
    END
  END GND
  PIN VDD
    ANTENNADIFFAREA 3.595900 ;
    PORT
      LAYER nwell ;
        RECT 16.380 10.160 17.220 10.170 ;
        RECT 19.380 10.160 20.220 10.170 ;
        RECT 16.380 8.580 22.820 10.160 ;
        RECT 16.380 7.610 22.840 8.580 ;
        RECT 16.610 7.600 22.840 7.610 ;
        RECT 19.420 7.590 22.840 7.600 ;
        RECT 11.630 6.570 12.490 6.700 ;
        RECT 9.070 4.960 12.490 6.570 ;
      LAYER li1 ;
        RECT 17.800 9.190 18.300 10.620 ;
        RECT 16.810 8.560 18.310 9.190 ;
        RECT 10.370 6.390 10.750 6.990 ;
        RECT 9.630 6.220 11.440 6.390 ;
        RECT 10.130 5.940 10.570 6.220 ;
        RECT 9.310 5.910 10.570 5.940 ;
        RECT 9.310 5.210 10.580 5.910 ;
      LAYER met1 ;
        RECT 17.800 10.660 18.280 10.720 ;
        RECT 10.610 10.580 18.280 10.660 ;
        RECT 10.450 10.340 18.280 10.580 ;
        RECT 10.450 8.790 10.720 10.340 ;
        RECT 17.800 10.310 18.280 10.340 ;
        RECT 10.400 6.600 10.760 8.790 ;
        RECT 9.510 6.470 12.180 6.600 ;
        RECT 9.510 6.190 12.210 6.470 ;
        RECT 9.510 5.960 12.180 6.190 ;
        RECT 9.510 5.950 9.680 5.960 ;
        RECT 10.130 5.950 12.180 5.960 ;
    END
  END VDD
  PIN a
    ANTENNAGATEAREA 0.607600 ;
    ANTENNADIFFAREA 0.726000 ;
    PORT
      LAYER li1 ;
        RECT 18.410 7.510 18.930 7.520 ;
        RECT 16.740 7.230 18.930 7.510 ;
        RECT 18.410 7.220 18.930 7.230 ;
        RECT 10.930 5.210 11.330 5.910 ;
        RECT 11.130 4.820 11.330 5.210 ;
        RECT 11.120 4.620 11.330 4.820 ;
        RECT 11.130 4.330 11.330 4.620 ;
        RECT 10.930 3.960 11.330 4.330 ;
      LAYER met1 ;
        RECT 16.730 7.480 17.150 7.520 ;
        RECT 18.580 7.480 18.910 7.500 ;
        RECT 13.480 7.300 18.910 7.480 ;
        RECT 13.480 7.230 13.980 7.300 ;
        RECT 11.050 4.800 11.390 4.850 ;
        RECT 13.530 4.800 13.830 7.230 ;
        RECT 16.730 7.220 17.150 7.300 ;
        RECT 18.580 7.270 18.910 7.300 ;
        RECT 11.050 4.630 13.830 4.800 ;
        RECT 11.050 4.570 11.360 4.630 ;
        RECT 11.130 4.560 11.360 4.570 ;
    END
  END a
  OBS
      LAYER li1 ;
        RECT 21.060 7.510 21.550 9.210 ;
        RECT 19.680 7.450 21.550 7.510 ;
        RECT 19.400 7.340 21.550 7.450 ;
        RECT 19.400 6.770 19.850 7.340 ;
        RECT 10.420 4.560 10.760 4.840 ;
  END
END nor
END LIBRARY

