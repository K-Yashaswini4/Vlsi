VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dlatch
  CLASS BLOCK ;
  FOREIGN dlatch ;
  ORIGIN 12.830 3.760 ;
  SIZE 27.680 BY 36.290 ;
  PIN D_in
    ANTENNADIFFAREA 2.111800 ;
    PORT
      LAYER li1 ;
        RECT 0.340 3.550 0.760 3.810 ;
        RECT 0.340 2.450 0.790 3.550 ;
        RECT 0.070 2.120 0.790 2.450 ;
        RECT 0.340 1.160 0.790 2.120 ;
        RECT 0.340 0.820 0.780 1.160 ;
      LAYER met1 ;
        RECT 0.310 2.920 0.770 2.930 ;
        RECT 0.130 2.580 0.770 2.920 ;
    END
  END D_in
  PIN clk_bar
    ANTENNAGATEAREA 0.928200 ;
    ANTENNADIFFAREA 0.726000 ;
    PORT
      LAYER li1 ;
        RECT -3.600 22.970 -2.910 23.460 ;
        RECT 1.590 23.430 2.170 23.520 ;
        RECT 1.590 23.020 2.180 23.430 ;
        RECT -3.450 22.560 -3.130 22.970 ;
        RECT 1.570 22.760 2.170 23.020 ;
        RECT -3.440 22.350 -3.130 22.560 ;
        RECT 1.560 22.500 2.060 22.760 ;
        RECT 1.560 22.350 2.680 22.500 ;
        RECT -3.440 22.330 -0.820 22.350 ;
        RECT -0.430 22.330 2.680 22.350 ;
        RECT -3.440 22.250 2.680 22.330 ;
        RECT -3.440 22.130 2.060 22.250 ;
        RECT -1.220 21.340 -0.940 22.130 ;
        RECT 1.220 5.720 1.830 5.730 ;
        RECT 1.220 5.710 3.790 5.720 ;
        RECT 4.510 5.710 6.290 5.720 ;
        RECT 1.220 5.440 6.800 5.710 ;
        RECT 0.110 5.310 6.800 5.440 ;
        RECT 0.110 5.300 4.280 5.310 ;
        RECT 4.510 5.300 6.800 5.310 ;
        RECT 0.110 5.070 1.830 5.300 ;
        RECT 3.810 5.290 4.280 5.300 ;
        RECT 1.050 4.880 1.830 5.070 ;
        RECT 1.070 4.730 1.830 4.880 ;
        RECT 6.290 4.800 6.800 5.300 ;
        RECT 1.070 4.690 1.780 4.730 ;
        RECT 1.090 4.260 1.780 4.690 ;
        RECT 6.280 4.290 6.870 4.800 ;
        RECT 6.280 4.200 6.860 4.290 ;
        RECT -6.110 2.280 -5.710 2.980 ;
        RECT -5.910 1.910 -5.710 2.280 ;
        RECT -5.910 1.490 -5.420 1.910 ;
        RECT -5.910 1.400 -5.710 1.490 ;
        RECT -6.110 1.030 -5.710 1.400 ;
      LAYER met1 ;
        RECT 2.060 22.620 2.510 22.710 ;
        RECT 2.060 22.440 3.390 22.620 ;
        RECT 2.060 22.230 3.420 22.440 ;
        RECT -1.260 21.740 -1.090 21.760 ;
        RECT 2.730 21.740 3.420 22.230 ;
        RECT -1.260 21.470 3.420 21.740 ;
        RECT -3.020 5.440 -2.530 5.460 ;
        RECT -3.020 5.060 1.300 5.440 ;
        RECT 2.730 5.360 3.420 21.470 ;
        RECT -3.020 5.010 1.660 5.060 ;
        RECT -3.020 4.870 1.670 5.010 ;
        RECT -3.020 4.840 1.210 4.870 ;
        RECT -3.020 1.870 -2.530 4.840 ;
        RECT 1.060 4.830 1.210 4.840 ;
        RECT 6.260 4.190 6.840 5.650 ;
        RECT -5.840 1.860 -2.530 1.870 ;
        RECT -5.840 1.540 -2.570 1.860 ;
    END
  END clk_bar
  PIN clock
    ANTENNAGATEAREA 1.109700 ;
    PORT
      LAYER li1 ;
        RECT 1.540 28.480 2.150 28.490 ;
        RECT -2.920 28.470 -1.140 28.480 ;
        RECT -0.420 28.470 2.150 28.480 ;
        RECT -3.430 28.200 2.150 28.470 ;
        RECT 14.170 28.220 14.380 28.260 ;
        RECT 3.180 28.200 14.380 28.220 ;
        RECT -3.430 28.140 14.380 28.200 ;
        RECT -3.430 28.070 14.450 28.140 ;
        RECT -3.430 28.060 -1.140 28.070 ;
        RECT -0.910 28.060 14.450 28.070 ;
        RECT -3.430 27.560 -2.920 28.060 ;
        RECT -0.910 28.050 -0.440 28.060 ;
        RECT 1.540 27.830 14.450 28.060 ;
        RECT -3.500 27.050 -2.910 27.560 ;
        RECT 1.540 27.510 2.150 27.830 ;
        RECT 3.180 27.740 14.450 27.830 ;
        RECT 1.540 27.490 2.280 27.510 ;
        RECT -3.490 26.960 -2.910 27.050 ;
        RECT 1.590 27.020 2.280 27.490 ;
        RECT 14.170 4.410 14.450 27.740 ;
        RECT 14.240 4.400 14.450 4.410 ;
        RECT -6.620 1.860 -6.280 1.910 ;
        RECT -7.300 1.630 -6.280 1.860 ;
        RECT -7.300 1.590 -6.620 1.630 ;
        RECT 1.200 0.670 1.780 0.760 ;
        RECT 1.190 0.260 1.780 0.670 ;
        RECT 1.200 0.000 1.800 0.260 ;
        RECT 6.280 0.210 6.970 0.700 ;
        RECT 1.310 -0.260 1.810 0.000 ;
        RECT 0.690 -0.410 1.810 -0.260 ;
        RECT 6.500 -0.200 6.820 0.210 ;
        RECT 4.210 -0.410 4.590 -0.290 ;
        RECT 6.500 -0.410 6.810 -0.200 ;
        RECT 0.690 -0.430 3.800 -0.410 ;
        RECT 4.190 -0.430 6.810 -0.410 ;
        RECT 0.690 -0.510 6.810 -0.430 ;
        RECT 1.310 -0.630 6.810 -0.510 ;
        RECT 14.240 -3.130 14.480 4.400 ;
        RECT 4.310 -3.600 14.480 -3.130 ;
        RECT 14.240 -3.620 14.480 -3.600 ;
      LAYER met1 ;
        RECT 2.070 27.840 2.700 28.200 ;
        RECT 2.070 27.740 2.610 27.840 ;
        RECT 1.700 27.600 2.610 27.740 ;
        RECT 1.700 27.060 2.070 27.600 ;
        RECT -8.790 1.580 -6.580 1.870 ;
        RECT -8.790 -0.050 -8.380 1.580 ;
        RECT -8.790 -0.130 -8.370 -0.050 ;
        RECT -3.680 -0.130 -0.090 -0.050 ;
        RECT -8.790 -0.140 -0.090 -0.130 ;
        RECT 0.860 -0.140 1.310 -0.050 ;
        RECT -8.790 -0.320 1.310 -0.140 ;
        RECT 0.550 -0.530 1.310 -0.320 ;
        RECT 4.250 -2.080 4.570 -0.320 ;
        RECT 4.250 -3.760 4.660 -2.080 ;
    END
  END clock
  PIN GND
    ANTENNADIFFAREA 2.260000 ;
    PORT
      LAYER li1 ;
        RECT -6.890 29.790 -5.640 30.160 ;
        RECT -7.850 28.970 -7.620 29.520 ;
        RECT -6.890 29.310 -6.440 29.790 ;
        RECT -8.470 28.720 -7.620 28.970 ;
        RECT -12.830 25.450 -8.210 25.930 ;
        RECT -12.830 4.930 -12.210 25.450 ;
        RECT -8.670 23.560 -8.470 23.570 ;
        RECT -8.670 23.090 -8.220 23.560 ;
        RECT -9.470 22.720 -8.220 23.090 ;
        RECT 9.010 7.030 10.260 7.400 ;
        RECT 0.670 6.710 1.780 6.800 ;
        RECT 8.320 6.720 9.170 6.730 ;
        RECT 7.980 6.710 9.170 6.720 ;
        RECT 0.670 6.550 9.170 6.710 ;
        RECT 9.810 6.550 10.260 7.030 ;
        RECT 0.670 6.490 8.490 6.550 ;
        RECT 0.670 6.320 1.780 6.490 ;
        RECT 7.730 6.220 8.020 6.490 ;
        RECT 7.730 6.210 8.190 6.220 ;
        RECT 10.990 6.210 11.220 6.760 ;
        RECT 7.730 6.050 11.840 6.210 ;
        RECT 7.740 5.970 11.840 6.050 ;
        RECT 10.990 5.960 11.840 5.970 ;
        RECT -12.760 0.820 -12.210 4.930 ;
        RECT -7.710 1.030 -6.460 1.400 ;
        RECT -6.910 0.820 -6.460 1.030 ;
        RECT -12.780 0.550 -6.460 0.820 ;
        RECT -4.310 1.110 -3.770 4.020 ;
        RECT -4.310 0.690 -3.880 1.110 ;
        RECT 11.420 0.810 11.840 3.160 ;
        RECT 11.420 0.800 12.040 0.810 ;
        RECT -12.780 0.470 -6.860 0.550 ;
        RECT -12.690 0.430 -6.860 0.470 ;
        RECT -12.690 0.420 -7.050 0.430 ;
        RECT -8.090 0.150 -7.780 0.420 ;
        RECT -8.040 0.100 -7.830 0.150 ;
        RECT -4.320 0.080 -3.880 0.690 ;
        RECT 11.590 0.330 12.040 0.800 ;
        RECT 11.590 -0.040 12.840 0.330 ;
      LAYER met1 ;
        RECT -6.890 29.790 -6.740 29.860 ;
        RECT -7.760 29.740 -5.740 29.790 ;
        RECT -7.920 29.610 -5.740 29.740 ;
        RECT -7.920 29.600 -5.980 29.610 ;
        RECT -7.900 29.190 -5.980 29.600 ;
        RECT -8.490 28.850 -7.970 29.020 ;
        RECT -8.650 28.720 -7.970 28.850 ;
        RECT -8.650 28.500 -8.210 28.720 ;
        RECT -8.600 23.720 -8.210 28.500 ;
        RECT -8.650 23.530 -8.230 23.720 ;
        RECT -8.650 23.230 -8.240 23.530 ;
        RECT -8.650 23.100 -8.220 23.230 ;
        RECT -8.560 23.090 -8.220 23.100 ;
        RECT -8.370 23.020 -8.220 23.090 ;
        RECT 10.110 7.030 10.260 7.100 ;
        RECT 9.110 6.990 11.300 7.030 ;
        RECT -4.020 6.870 0.990 6.880 ;
        RECT -4.020 6.860 1.070 6.870 ;
        RECT -4.020 6.670 1.100 6.860 ;
        RECT 9.110 6.850 11.350 6.990 ;
        RECT 9.110 6.760 11.860 6.850 ;
        RECT -4.370 6.250 1.100 6.670 ;
        RECT 7.750 6.430 11.860 6.760 ;
        RECT 7.750 6.410 9.340 6.430 ;
        RECT 11.300 6.290 11.860 6.430 ;
        RECT -4.370 6.240 1.070 6.250 ;
        RECT -4.370 4.020 -3.780 6.240 ;
        RECT -4.370 3.620 -3.700 4.020 ;
        RECT -6.610 1.030 -6.460 1.100 ;
        RECT -7.610 1.010 -5.000 1.030 ;
        RECT -7.610 0.740 -3.880 1.010 ;
        RECT 11.340 0.930 11.860 6.290 ;
        RECT -7.610 0.430 -5.420 0.740 ;
        RECT -5.060 0.620 -3.880 0.740 ;
        RECT -8.110 0.270 -7.760 0.360 ;
        RECT -4.320 0.270 -3.880 0.620 ;
        RECT 10.550 0.330 12.740 0.930 ;
        RECT -8.110 0.190 -3.920 0.270 ;
        RECT 11.590 0.260 11.740 0.330 ;
        RECT -8.100 0.050 -3.920 0.190 ;
    END
  END GND
  PIN VDD
    ANTENNADIFFAREA 6.835500 ;
    PORT
      LAYER nwell ;
        RECT -8.800 32.400 -7.940 32.530 ;
        RECT -8.800 30.790 -5.380 32.400 ;
        RECT -9.730 20.480 -6.310 22.090 ;
        RECT -7.170 20.350 -6.310 20.480 ;
        RECT 11.310 9.640 12.170 9.770 ;
        RECT 8.750 8.030 12.170 9.640 ;
        RECT -5.410 3.640 -4.550 3.770 ;
        RECT -7.970 2.030 -4.550 3.640 ;
        RECT 9.680 -2.280 13.100 -0.670 ;
        RECT 9.680 -2.410 10.540 -2.280 ;
      LAYER li1 ;
        RECT -7.750 32.050 -5.980 32.220 ;
        RECT -6.880 31.770 -6.440 32.050 ;
        RECT -6.880 31.740 -5.620 31.770 ;
        RECT -6.890 31.040 -5.620 31.740 ;
        RECT -9.490 21.140 -8.220 21.840 ;
        RECT -9.490 21.110 -8.230 21.140 ;
        RECT -8.670 20.830 -8.230 21.110 ;
        RECT -9.130 20.660 -7.360 20.830 ;
        RECT -5.660 9.600 9.350 9.670 ;
        RECT -6.440 9.460 9.350 9.600 ;
        RECT -6.440 9.290 11.120 9.460 ;
        RECT -6.440 9.210 10.250 9.290 ;
        RECT -6.440 8.940 -5.670 9.210 ;
        RECT 9.810 9.010 10.250 9.210 ;
        RECT 8.990 8.980 10.250 9.010 ;
        RECT 8.990 8.280 10.260 8.980 ;
        RECT -7.370 3.290 -5.600 3.460 ;
        RECT -6.910 3.010 -6.470 3.290 ;
        RECT -7.730 2.980 -6.470 3.010 ;
        RECT -7.730 2.280 -6.460 2.980 ;
        RECT 11.590 -1.620 12.860 -0.920 ;
        RECT 11.600 -1.650 12.860 -1.620 ;
        RECT 11.600 -1.930 12.040 -1.650 ;
        RECT 10.730 -2.100 12.500 -1.930 ;
      LAYER met1 ;
        RECT -10.450 32.420 -5.820 32.430 ;
        RECT -10.450 31.930 -5.790 32.420 ;
        RECT -10.450 31.910 -5.820 31.930 ;
        RECT -10.450 31.900 -10.240 31.910 ;
        RECT -10.450 21.060 -10.260 31.900 ;
        RECT -8.490 31.790 -5.820 31.910 ;
        RECT -8.490 31.780 -6.440 31.790 ;
        RECT -5.990 31.780 -5.820 31.790 ;
        RECT -10.820 21.040 -10.260 21.060 ;
        RECT -9.290 21.090 -9.120 21.100 ;
        RECT -8.670 21.090 -6.620 21.100 ;
        RECT -9.290 21.060 -6.620 21.090 ;
        RECT -9.290 21.040 -5.920 21.060 ;
        RECT -11.480 20.700 -5.920 21.040 ;
        RECT -11.480 20.520 -5.790 20.700 ;
        RECT -9.290 20.450 -5.790 20.520 ;
        RECT -6.860 20.330 -5.790 20.450 ;
        RECT -6.470 9.210 -5.790 20.330 ;
        RECT 8.860 10.100 9.200 10.110 ;
        RECT 8.860 10.070 12.500 10.100 ;
        RECT 8.860 9.900 12.850 10.070 ;
        RECT 8.860 9.670 9.200 9.900 ;
        RECT 8.860 9.540 11.860 9.670 ;
        RECT 8.860 9.260 11.890 9.540 ;
        RECT 12.490 9.350 12.850 9.900 ;
        RECT -6.470 9.020 -5.690 9.210 ;
        RECT 8.860 9.070 11.860 9.260 ;
        RECT 12.490 9.180 13.820 9.350 ;
        RECT 12.820 9.120 13.820 9.180 ;
        RECT 9.190 9.030 11.860 9.070 ;
        RECT 9.190 9.020 9.360 9.030 ;
        RECT 9.810 9.020 11.860 9.030 ;
        RECT -6.450 6.100 -5.690 9.020 ;
        RECT -6.440 3.670 -5.710 6.100 ;
        RECT -7.530 3.540 -4.860 3.670 ;
        RECT -7.530 3.260 -4.830 3.540 ;
        RECT -7.530 3.030 -4.860 3.260 ;
        RECT -7.530 3.020 -7.360 3.030 ;
        RECT -6.910 3.020 -4.860 3.030 ;
        RECT 9.990 -1.670 12.040 -1.660 ;
        RECT 12.490 -1.670 12.660 -1.660 ;
        RECT 9.990 -1.700 12.660 -1.670 ;
        RECT 9.730 -1.720 12.660 -1.700 ;
        RECT 13.630 -1.700 13.820 9.120 ;
        RECT 13.630 -1.720 14.190 -1.700 ;
        RECT 9.730 -2.240 14.850 -1.720 ;
        RECT 9.730 -2.310 12.660 -2.240 ;
        RECT 9.730 -2.340 9.990 -2.310 ;
    END
  END VDD
  PIN Q1
    ANTENNAGATEAREA 0.181500 ;
    ANTENNADIFFAREA 2.265600 ;
    PORT
      LAYER li1 ;
        RECT 8.800 7.630 10.440 7.910 ;
        RECT 5.500 3.690 5.940 3.730 ;
        RECT 2.120 2.460 2.570 3.600 ;
        RECT 5.490 2.830 5.940 3.690 ;
        RECT 5.230 2.500 5.940 2.830 ;
        RECT 5.210 2.460 5.970 2.500 ;
        RECT 2.120 2.170 2.880 2.460 ;
        RECT 4.510 2.180 5.970 2.460 ;
        RECT 4.580 2.170 5.970 2.180 ;
        RECT 2.120 2.130 2.830 2.170 ;
        RECT 2.120 1.270 2.570 2.130 ;
        RECT 5.490 1.360 5.940 2.170 ;
        RECT 2.120 1.230 2.560 1.270 ;
      LAYER met1 ;
        RECT 8.610 7.800 9.100 7.910 ;
        RECT 4.200 7.670 9.100 7.800 ;
        RECT 4.200 7.640 8.790 7.670 ;
        RECT 4.200 6.950 4.500 7.640 ;
        RECT 4.220 6.370 4.490 6.950 ;
        RECT 4.200 5.710 4.500 6.370 ;
        RECT 2.390 2.460 2.880 2.490 ;
        RECT 4.280 2.460 4.510 5.710 ;
        RECT 5.220 2.500 5.950 2.510 ;
        RECT 5.210 2.460 5.960 2.500 ;
        RECT 2.390 2.180 5.960 2.460 ;
        RECT 2.390 2.170 4.280 2.180 ;
        RECT 2.420 2.140 2.780 2.170 ;
        RECT 4.590 2.150 5.960 2.180 ;
    END
  END Q1
  PIN Q1out
    ANTENNAGATEAREA 0.181500 ;
    ANTENNADIFFAREA 2.837800 ;
    PORT
      LAYER li1 ;
        RECT 2.610 26.310 3.030 26.570 ;
        RECT 2.580 25.210 3.030 26.310 ;
        RECT 2.580 24.880 3.300 25.210 ;
        RECT 2.580 23.920 3.030 24.880 ;
        RECT 2.590 23.580 3.030 23.920 ;
        RECT 10.610 8.280 11.010 8.980 ;
        RECT 10.810 7.920 11.010 8.280 ;
        RECT 12.990 7.920 13.440 10.140 ;
        RECT 10.810 7.630 13.450 7.920 ;
        RECT 10.810 7.400 11.010 7.630 ;
        RECT 13.090 7.620 13.450 7.630 ;
        RECT 10.610 7.030 11.010 7.400 ;
        RECT 11.410 -0.290 11.750 -0.270 ;
        RECT 11.410 -0.550 13.460 -0.290 ;
        RECT 11.740 -0.560 13.460 -0.550 ;
      LAYER met1 ;
        RECT 2.600 25.680 3.060 25.690 ;
        RECT 2.600 25.670 3.240 25.680 ;
        RECT 2.600 25.660 3.410 25.670 ;
        RECT 2.600 25.440 13.450 25.660 ;
        RECT 2.600 25.350 3.410 25.440 ;
        RECT 2.600 25.340 3.240 25.350 ;
        RECT 11.980 25.220 13.450 25.440 ;
        RECT 13.080 13.450 13.410 25.220 ;
        RECT 13.150 12.580 13.410 13.450 ;
        RECT 13.150 12.270 13.500 12.580 ;
        RECT 13.150 11.640 13.450 12.270 ;
        RECT 13.000 9.810 13.450 11.640 ;
        RECT 13.100 7.620 13.440 7.900 ;
        RECT 13.090 -0.530 13.480 7.620 ;
        RECT 13.090 -0.550 13.470 -0.530 ;
    END
  END Q1out
  PIN Q1bar_out
    ANTENNADIFFAREA 1.986900 ;
    PORT
      LAYER li1 ;
        RECT 7.280 3.800 7.720 4.140 ;
        RECT 7.270 2.840 7.720 3.800 ;
        RECT 7.270 2.510 8.950 2.840 ;
        RECT 7.270 1.410 7.720 2.510 ;
        RECT 7.980 2.450 8.950 2.510 ;
        RECT 7.300 1.150 7.720 1.410 ;
        RECT 10.840 -0.040 11.240 0.330 ;
        RECT 10.840 -0.200 11.040 -0.040 ;
        RECT 9.000 -0.510 11.040 -0.200 ;
        RECT 10.840 -0.920 11.040 -0.510 ;
        RECT 10.840 -1.620 11.240 -0.920 ;
      LAYER met1 ;
        RECT 7.860 -0.180 8.950 2.840 ;
        RECT 7.860 -0.630 9.300 -0.180 ;
    END
  END Q1bar_out
  PIN Q1out_bar
    ANTENNAGATEAREA 0.181500 ;
    ANTENNADIFFAREA 2.265600 ;
    PORT
      LAYER li1 ;
        RECT -7.070 30.390 -5.430 30.670 ;
        RECT -2.570 26.450 -2.130 26.490 ;
        RECT -2.570 25.590 -2.120 26.450 ;
        RECT -2.570 25.260 -1.860 25.590 ;
        RECT -2.600 25.220 -1.840 25.260 ;
        RECT 0.800 25.220 1.250 26.360 ;
        RECT -2.600 24.940 -1.140 25.220 ;
        RECT -2.600 24.930 -1.210 24.940 ;
        RECT 0.490 24.930 1.250 25.220 ;
        RECT -2.570 24.120 -2.120 24.930 ;
        RECT 0.540 24.890 1.250 24.930 ;
        RECT 0.800 24.030 1.250 24.890 ;
        RECT 0.810 23.990 1.250 24.030 ;
      LAYER met1 ;
        RECT -5.730 30.560 -5.240 30.670 ;
        RECT -5.730 30.430 -0.830 30.560 ;
        RECT -5.420 30.400 -0.830 30.430 ;
        RECT -1.130 29.710 -0.830 30.400 ;
        RECT -1.120 29.130 -0.850 29.710 ;
        RECT -1.130 28.470 -0.830 29.130 ;
        RECT -2.580 25.260 -1.850 25.270 ;
        RECT -2.590 25.220 -1.840 25.260 ;
        RECT -1.140 25.220 -0.910 28.470 ;
        RECT 0.490 25.220 0.980 25.250 ;
        RECT -2.590 24.940 0.980 25.220 ;
        RECT -2.590 24.910 -1.220 24.940 ;
        RECT -0.910 24.930 0.980 24.940 ;
        RECT 0.590 24.900 0.950 24.930 ;
    END
  END Q1out_bar
  PIN Q2
    ANTENNAGATEAREA 0.181500 ;
    ANTENNADIFFAREA 0.726000 ;
    PORT
      LAYER li1 ;
        RECT -7.640 31.040 -7.240 31.740 ;
        RECT -7.640 30.680 -7.440 31.040 ;
        RECT -10.080 30.390 -7.440 30.680 ;
        RECT -10.080 30.380 -9.720 30.390 ;
        RECT -7.640 30.160 -7.440 30.390 ;
        RECT -7.640 29.790 -7.240 30.160 ;
        RECT -8.380 22.470 -8.040 22.490 ;
        RECT -10.090 22.210 -8.040 22.470 ;
        RECT -10.090 22.200 -8.370 22.210 ;
      LAYER met1 ;
        RECT -10.070 30.380 -9.730 30.660 ;
        RECT -10.110 22.230 -9.720 30.380 ;
        RECT -10.100 22.210 -9.720 22.230 ;
    END
  END Q2
  OBS
      LAYER nwell ;
        RECT -4.700 27.730 -3.850 27.760 ;
        RECT -4.700 27.720 -3.760 27.730 ;
        RECT -4.700 26.900 -1.810 27.720 ;
        RECT -4.690 25.880 -1.810 26.900 ;
        RECT -4.670 25.260 -1.810 25.880 ;
        RECT 0.490 22.840 5.100 25.220 ;
        RECT 0.490 22.760 3.380 22.840 ;
        RECT 2.440 22.750 3.380 22.760 ;
        RECT 2.530 22.720 3.380 22.750 ;
        RECT 7.220 4.970 8.070 5.000 ;
        RECT 7.130 4.960 8.070 4.970 ;
        RECT 5.180 4.140 8.070 4.960 ;
        RECT 5.180 3.120 8.060 4.140 ;
        RECT 5.180 2.500 8.040 3.120 ;
        RECT -1.730 0.080 2.880 2.460 ;
        RECT -0.010 0.000 2.880 0.080 ;
        RECT -0.010 -0.010 0.930 0.000 ;
        RECT -0.010 -0.040 0.840 -0.010 ;
      LAYER li1 ;
        RECT -4.350 26.560 -3.910 26.900 ;
        RECT -4.350 25.600 -3.900 26.560 ;
        RECT -5.580 25.270 -3.900 25.600 ;
        RECT -5.580 25.210 -4.610 25.270 ;
        RECT -4.350 24.170 -3.900 25.270 ;
        RECT -4.350 23.910 -3.930 24.170 ;
        RECT -7.870 22.720 -7.470 23.090 ;
        RECT -7.670 22.560 -7.470 22.720 ;
        RECT -7.670 22.250 -5.630 22.560 ;
        RECT -7.670 21.840 -7.470 22.250 ;
        RECT -7.870 21.140 -7.470 21.840 ;
      LAYER met1 ;
        RECT -5.580 22.580 -4.490 25.600 ;
        RECT -5.930 22.130 -4.490 22.580 ;
  END
END dlatch
END LIBRARY

